module IBUF (
    input  wire logic I,
    output      logic O
    );

    // NULL MODULE

endmodule