module MMCME2_ADV #(
    parameter BANDWIDTH = "OPTIMIZED",
    parameter CLKFBOUT_MULT_F = 5.000,
    parameter CLKFBOUT_PHASE = 0.000,
    parameter CLKFBOUT_USE_FINE_PS = "FALSE",
    parameter CLKIN1_PERIOD = 0.000,
    parameter CLKIN2_PERIOD = 0.000,
    parameter CLKOUT0_DIVIDE_F = 1.000,
    parameter CLKOUT0_DUTY_CYCLE = 0.500,
    parameter CLKOUT0_PHASE = 0.000,
    parameter CLKOUT0_USE_FINE_PS = "FALSE",
    parameter CLKOUT1_DIVIDE = 1,
    parameter CLKOUT1_DUTY_CYCLE = 0.500,
    parameter CLKOUT1_PHASE = 0.000,
    parameter CLKOUT1_USE_FINE_PS = "FALSE",
    parameter CLKOUT2_DIVIDE = 1,
    parameter CLKOUT2_DUTY_CYCLE = 0.500,
    parameter CLKOUT2_PHASE = 0.000,
    parameter CLKOUT2_USE_FINE_PS = "FALSE",
    parameter CLKOUT3_DIVIDE = 1,
    parameter CLKOUT3_DUTY_CYCLE = 0.500,
    parameter CLKOUT3_PHASE = 0.000,
    parameter CLKOUT3_USE_FINE_PS = "FALSE",
    parameter CLKOUT4_CASCADE = "FALSE",
    parameter CLKOUT4_DIVIDE = 1,
    parameter CLKOUT4_DUTY_CYCLE = 0.500,
    parameter CLKOUT4_PHASE = 0.000,
    parameter CLKOUT4_USE_FINE_PS = "FALSE",
    parameter CLKOUT5_DIVIDE = 1,
    parameter CLKOUT5_DUTY_CYCLE = 0.500,
    parameter CLKOUT5_PHASE = 0.000,
    parameter CLKOUT5_USE_FINE_PS = "FALSE",
    parameter CLKOUT6_DIVIDE = 1,
    parameter CLKOUT6_DUTY_CYCLE = 0.500,
    parameter CLKOUT6_PHASE = 0.000,
    parameter CLKOUT6_USE_FINE_PS = "FALSE",
    parameter COMPENSATION = "ZHOLD",
    parameter DIVCLK_DIVIDE = 1,
    parameter REF_JITTER1 = 0.0,
    parameter REF_JITTER2 = 0.0,
    parameter SS_EN = "FALSE",
    parameter SS_MODE = "CENTER_HIGH",
    parameter SS_MOD_PERIOD = 10000,
    parameter STARTUP_WAIT = "FALSE"
)(
    output logic CLKFBOUT,
    output logic CLKFBOUTB,
    output logic CLKFBSTOPPED,
    output logic CLKINSTOPPED,
    output logic CLKOUT0,
    output logic CLKOUT0B,
    output logic CLKOUT1,
    output logic CLKOUT1B,
    output logic CLKOUT2,
    output logic CLKOUT2B,
    output logic CLKOUT3,
    output logic CLKOUT3B,
    output logic CLKOUT4,
    output logic CLKOUT5,
    output logic CLKOUT6,
    output logic [15:0] DO,
    output logic DRDY,
    output logic LOCKED,
    output logic PSDONE,

    input wire CLKFBIN,
    input wire CLKIN1,
    input wire CLKIN2,
    input wire CLKINSEL,
    input wire [6:0] DADDR,
    input wire DCLK,
    input wire DEN,
    input wire [15:0] DI,
    input wire DWE,
    input wire PSCLK,
    input wire PSEN,
    input wire PSINCDEC,
    input wire PWRDWN,
    input wire RST
);


endmodule